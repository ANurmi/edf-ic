module seq_prio_queue #()();

endmodule : seq_prio_queue
