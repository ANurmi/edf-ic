module seq_prio_queue #()(
  input logic clk_i,
  input logic rst_ni
);

endmodule : seq_prio_queue
