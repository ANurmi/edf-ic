module edf_ic #(
  parameter int unsigned SerLatency = 1
)(
  input  logic                   clk_i,
  input  logic                   rst_ni,
  output logic                   irq_id_o
);

endmodule : edf_ic
