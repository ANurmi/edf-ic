module gateway_cell #()();
endmodule : gateway_cell
