module tb_edf_intctl_top #(
)();

endmodule : tb_edf_intctl_top
